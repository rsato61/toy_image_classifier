library verilog;
use verilog.vl_types.all;
entity freds_house_testbench is
end freds_house_testbench;
