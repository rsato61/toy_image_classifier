library verilog;
use verilog.vl_types.all;
entity seg2x7_testbench is
end seg2x7_testbench;
