library verilog;
use verilog.vl_types.all;
entity victory_testbench is
end victory_testbench;
