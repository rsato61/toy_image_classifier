// cpu.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module cpu (
		input  wire [7:0]  classification_pio_export, // classification_pio.export
		input  wire        clk_clk,                   //                clk.clk
		input  wire [31:0] distance_pio_export,       //       distance_pio.export
		output wire [7:0]  done_read_pio_export,      //      done_read_pio.export
		input  wire [7:0]  read_diff_pio_export,      //      read_diff_pio.export
		input  wire        reset_reset_n,             //              reset.reset_n
		output wire        sdram_clk_clk              //          sdram_clk.clk
	);

	wire         sys_sdram_pll_0_sys_clk_clk;                            // sys_sdram_pll_0:sys_clk_clk -> [cpu_nios:clk, irq_mapper:clk, jtag:clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, onchip_memory:clk, rst_controller_001:clk, rst_controller_002:clk, sysid_qsys_0:clock]
	wire  [31:0] cpu_nios_data_master_readdata;                          // mm_interconnect_0:cpu_nios_data_master_readdata -> cpu_nios:d_readdata
	wire         cpu_nios_data_master_waitrequest;                       // mm_interconnect_0:cpu_nios_data_master_waitrequest -> cpu_nios:d_waitrequest
	wire         cpu_nios_data_master_debugaccess;                       // cpu_nios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_nios_data_master_debugaccess
	wire  [17:0] cpu_nios_data_master_address;                           // cpu_nios:d_address -> mm_interconnect_0:cpu_nios_data_master_address
	wire   [3:0] cpu_nios_data_master_byteenable;                        // cpu_nios:d_byteenable -> mm_interconnect_0:cpu_nios_data_master_byteenable
	wire         cpu_nios_data_master_read;                              // cpu_nios:d_read -> mm_interconnect_0:cpu_nios_data_master_read
	wire         cpu_nios_data_master_write;                             // cpu_nios:d_write -> mm_interconnect_0:cpu_nios_data_master_write
	wire  [31:0] cpu_nios_data_master_writedata;                         // cpu_nios:d_writedata -> mm_interconnect_0:cpu_nios_data_master_writedata
	wire  [31:0] cpu_nios_instruction_master_readdata;                   // mm_interconnect_0:cpu_nios_instruction_master_readdata -> cpu_nios:i_readdata
	wire         cpu_nios_instruction_master_waitrequest;                // mm_interconnect_0:cpu_nios_instruction_master_waitrequest -> cpu_nios:i_waitrequest
	wire  [17:0] cpu_nios_instruction_master_address;                    // cpu_nios:i_address -> mm_interconnect_0:cpu_nios_instruction_master_address
	wire         cpu_nios_instruction_master_read;                       // cpu_nios:i_read -> mm_interconnect_0:cpu_nios_instruction_master_read
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;    // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;      // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;   // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;       // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;          // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;         // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;     // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;  // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;   // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_cpu_nios_debug_mem_slave_readdata;    // cpu_nios:debug_mem_slave_readdata -> mm_interconnect_0:cpu_nios_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_nios_debug_mem_slave_waitrequest; // cpu_nios:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_nios_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_nios_debug_mem_slave_debugaccess; // mm_interconnect_0:cpu_nios_debug_mem_slave_debugaccess -> cpu_nios:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_nios_debug_mem_slave_address;     // mm_interconnect_0:cpu_nios_debug_mem_slave_address -> cpu_nios:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_nios_debug_mem_slave_read;        // mm_interconnect_0:cpu_nios_debug_mem_slave_read -> cpu_nios:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_nios_debug_mem_slave_byteenable;  // mm_interconnect_0:cpu_nios_debug_mem_slave_byteenable -> cpu_nios:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_nios_debug_mem_slave_write;       // mm_interconnect_0:cpu_nios_debug_mem_slave_write -> cpu_nios:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_nios_debug_mem_slave_writedata;   // mm_interconnect_0:cpu_nios_debug_mem_slave_writedata -> cpu_nios:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;          // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;            // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory_s1_address;             // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;          // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;               // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;           // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;               // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire  [31:0] mm_interconnect_0_classification_pio_s1_readdata;       // classification_pio:readdata -> mm_interconnect_0:classification_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_classification_pio_s1_address;        // mm_interconnect_0:classification_pio_s1_address -> classification_pio:address
	wire         mm_interconnect_0_done_read_pio_s1_chipselect;          // mm_interconnect_0:done_read_pio_s1_chipselect -> done_read_pio:chipselect
	wire  [31:0] mm_interconnect_0_done_read_pio_s1_readdata;            // done_read_pio:readdata -> mm_interconnect_0:done_read_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_done_read_pio_s1_address;             // mm_interconnect_0:done_read_pio_s1_address -> done_read_pio:address
	wire         mm_interconnect_0_done_read_pio_s1_write;               // mm_interconnect_0:done_read_pio_s1_write -> done_read_pio:write_n
	wire  [31:0] mm_interconnect_0_done_read_pio_s1_writedata;           // mm_interconnect_0:done_read_pio_s1_writedata -> done_read_pio:writedata
	wire  [31:0] mm_interconnect_0_read_diff_pio_s1_readdata;            // read_diff_pio:readdata -> mm_interconnect_0:read_diff_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_read_diff_pio_s1_address;             // mm_interconnect_0:read_diff_pio_s1_address -> read_diff_pio:address
	wire  [31:0] mm_interconnect_0_distance_pio_s1_readdata;             // distance_pio:readdata -> mm_interconnect_0:distance_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_distance_pio_s1_address;              // mm_interconnect_0:distance_pio_s1_address -> distance_pio:address
	wire         irq_mapper_receiver0_irq;                               // jtag:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] cpu_nios_irq_irq;                                       // irq_mapper:sender_irq -> cpu_nios:irq
	wire         rst_controller_reset_out_reset;                         // rst_controller:reset_out -> [classification_pio:reset_n, distance_pio:reset_n, done_read_pio:reset_n, mm_interconnect_0:classification_pio_reset_reset_bridge_in_reset_reset, read_diff_pio:reset_n]
	wire         cpu_nios_debug_reset_request_reset;                     // cpu_nios:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_003:reset_in1]
	wire         rst_controller_001_reset_out_reset;                     // rst_controller_001:reset_out -> [cpu_nios:reset_n, irq_mapper:reset, mm_interconnect_0:cpu_nios_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_translator:in_reset, sysid_qsys_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                 // rst_controller_001:reset_req -> [cpu_nios:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                     // rst_controller_002:reset_out -> [jtag:rst_n, mm_interconnect_0:jtag_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_003_reset_out_reset;                     // rst_controller_003:reset_out -> sys_sdram_pll_0:ref_reset_reset

	cpu_classification_pio classification_pio (
		.clk      (clk_clk),                                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address  (mm_interconnect_0_classification_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_classification_pio_s1_readdata), //                    .readdata
		.in_port  (classification_pio_export)                         // external_connection.export
	);

	cpu_cpu_nios cpu_nios (
		.clk                                 (sys_sdram_pll_0_sys_clk_clk),                            //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (cpu_nios_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_nios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_nios_data_master_read),                              //                          .read
		.d_readdata                          (cpu_nios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_nios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_nios_data_master_write),                             //                          .write
		.d_writedata                         (cpu_nios_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_nios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_nios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_nios_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_nios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_nios_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_nios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_nios_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_nios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_nios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_nios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_nios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_nios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_nios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_nios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_nios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                        // custom_instruction_master.readra
	);

	cpu_distance_pio distance_pio (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_distance_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_distance_pio_s1_readdata), //                    .readdata
		.in_port  (distance_pio_export)                         // external_connection.export
	);

	cpu_done_read_pio done_read_pio (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_done_read_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_done_read_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_done_read_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_done_read_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_done_read_pio_s1_readdata),   //                    .readdata
		.out_port   (done_read_pio_export)                           // external_connection.export
	);

	cpu_jtag jtag (
		.clk            (sys_sdram_pll_0_sys_clk_clk),                          //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                  //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	cpu_onchip_memory onchip_memory (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                   //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),        //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	cpu_classification_pio read_diff_pio (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_read_diff_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_read_diff_pio_s1_readdata), //                    .readdata
		.in_port  (read_diff_pio_export)                         // external_connection.export
	);

	cpu_sys_sdram_pll_0 sys_sdram_pll_0 (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_003_reset_out_reset), //    ref_reset.reset
		.sys_clk_clk        (sys_sdram_pll_0_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                      //    sdram_clk.clk
		.reset_source_reset ()                                    // reset_source.reset
	);

	cpu_sysid_qsys_0 sysid_qsys_0 (
		.clock    (sys_sdram_pll_0_sys_clk_clk),                           //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	cpu_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                        (clk_clk),                                                //                                      clk_0_clk.clk
		.sys_sdram_pll_0_sys_clk_clk                          (sys_sdram_pll_0_sys_clk_clk),                            //                        sys_sdram_pll_0_sys_clk.clk
		.classification_pio_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                         // classification_pio_reset_reset_bridge_in_reset.reset
		.cpu_nios_reset_reset_bridge_in_reset_reset           (rst_controller_001_reset_out_reset),                     //           cpu_nios_reset_reset_bridge_in_reset.reset
		.jtag_reset_reset_bridge_in_reset_reset               (rst_controller_002_reset_out_reset),                     //               jtag_reset_reset_bridge_in_reset.reset
		.cpu_nios_data_master_address                         (cpu_nios_data_master_address),                           //                           cpu_nios_data_master.address
		.cpu_nios_data_master_waitrequest                     (cpu_nios_data_master_waitrequest),                       //                                               .waitrequest
		.cpu_nios_data_master_byteenable                      (cpu_nios_data_master_byteenable),                        //                                               .byteenable
		.cpu_nios_data_master_read                            (cpu_nios_data_master_read),                              //                                               .read
		.cpu_nios_data_master_readdata                        (cpu_nios_data_master_readdata),                          //                                               .readdata
		.cpu_nios_data_master_write                           (cpu_nios_data_master_write),                             //                                               .write
		.cpu_nios_data_master_writedata                       (cpu_nios_data_master_writedata),                         //                                               .writedata
		.cpu_nios_data_master_debugaccess                     (cpu_nios_data_master_debugaccess),                       //                                               .debugaccess
		.cpu_nios_instruction_master_address                  (cpu_nios_instruction_master_address),                    //                    cpu_nios_instruction_master.address
		.cpu_nios_instruction_master_waitrequest              (cpu_nios_instruction_master_waitrequest),                //                                               .waitrequest
		.cpu_nios_instruction_master_read                     (cpu_nios_instruction_master_read),                       //                                               .read
		.cpu_nios_instruction_master_readdata                 (cpu_nios_instruction_master_readdata),                   //                                               .readdata
		.classification_pio_s1_address                        (mm_interconnect_0_classification_pio_s1_address),        //                          classification_pio_s1.address
		.classification_pio_s1_readdata                       (mm_interconnect_0_classification_pio_s1_readdata),       //                                               .readdata
		.cpu_nios_debug_mem_slave_address                     (mm_interconnect_0_cpu_nios_debug_mem_slave_address),     //                       cpu_nios_debug_mem_slave.address
		.cpu_nios_debug_mem_slave_write                       (mm_interconnect_0_cpu_nios_debug_mem_slave_write),       //                                               .write
		.cpu_nios_debug_mem_slave_read                        (mm_interconnect_0_cpu_nios_debug_mem_slave_read),        //                                               .read
		.cpu_nios_debug_mem_slave_readdata                    (mm_interconnect_0_cpu_nios_debug_mem_slave_readdata),    //                                               .readdata
		.cpu_nios_debug_mem_slave_writedata                   (mm_interconnect_0_cpu_nios_debug_mem_slave_writedata),   //                                               .writedata
		.cpu_nios_debug_mem_slave_byteenable                  (mm_interconnect_0_cpu_nios_debug_mem_slave_byteenable),  //                                               .byteenable
		.cpu_nios_debug_mem_slave_waitrequest                 (mm_interconnect_0_cpu_nios_debug_mem_slave_waitrequest), //                                               .waitrequest
		.cpu_nios_debug_mem_slave_debugaccess                 (mm_interconnect_0_cpu_nios_debug_mem_slave_debugaccess), //                                               .debugaccess
		.distance_pio_s1_address                              (mm_interconnect_0_distance_pio_s1_address),              //                                distance_pio_s1.address
		.distance_pio_s1_readdata                             (mm_interconnect_0_distance_pio_s1_readdata),             //                                               .readdata
		.done_read_pio_s1_address                             (mm_interconnect_0_done_read_pio_s1_address),             //                               done_read_pio_s1.address
		.done_read_pio_s1_write                               (mm_interconnect_0_done_read_pio_s1_write),               //                                               .write
		.done_read_pio_s1_readdata                            (mm_interconnect_0_done_read_pio_s1_readdata),            //                                               .readdata
		.done_read_pio_s1_writedata                           (mm_interconnect_0_done_read_pio_s1_writedata),           //                                               .writedata
		.done_read_pio_s1_chipselect                          (mm_interconnect_0_done_read_pio_s1_chipselect),          //                                               .chipselect
		.jtag_avalon_jtag_slave_address                       (mm_interconnect_0_jtag_avalon_jtag_slave_address),       //                         jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write                         (mm_interconnect_0_jtag_avalon_jtag_slave_write),         //                                               .write
		.jtag_avalon_jtag_slave_read                          (mm_interconnect_0_jtag_avalon_jtag_slave_read),          //                                               .read
		.jtag_avalon_jtag_slave_readdata                      (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),      //                                               .readdata
		.jtag_avalon_jtag_slave_writedata                     (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),     //                                               .writedata
		.jtag_avalon_jtag_slave_waitrequest                   (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),   //                                               .waitrequest
		.jtag_avalon_jtag_slave_chipselect                    (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),    //                                               .chipselect
		.onchip_memory_s1_address                             (mm_interconnect_0_onchip_memory_s1_address),             //                               onchip_memory_s1.address
		.onchip_memory_s1_write                               (mm_interconnect_0_onchip_memory_s1_write),               //                                               .write
		.onchip_memory_s1_readdata                            (mm_interconnect_0_onchip_memory_s1_readdata),            //                                               .readdata
		.onchip_memory_s1_writedata                           (mm_interconnect_0_onchip_memory_s1_writedata),           //                                               .writedata
		.onchip_memory_s1_byteenable                          (mm_interconnect_0_onchip_memory_s1_byteenable),          //                                               .byteenable
		.onchip_memory_s1_chipselect                          (mm_interconnect_0_onchip_memory_s1_chipselect),          //                                               .chipselect
		.onchip_memory_s1_clken                               (mm_interconnect_0_onchip_memory_s1_clken),               //                                               .clken
		.read_diff_pio_s1_address                             (mm_interconnect_0_read_diff_pio_s1_address),             //                               read_diff_pio_s1.address
		.read_diff_pio_s1_readdata                            (mm_interconnect_0_read_diff_pio_s1_readdata),            //                                               .readdata
		.sysid_qsys_0_control_slave_address                   (mm_interconnect_0_sysid_qsys_0_control_slave_address),   //                     sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                  (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)   //                                               .readdata
	);

	cpu_irq_mapper irq_mapper (
		.clk           (sys_sdram_pll_0_sys_clk_clk),        //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (cpu_nios_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_nios_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_nios_debug_reset_request_reset),     // reset_in1.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),        //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_nios_debug_reset_request_reset), // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
